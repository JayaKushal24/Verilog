`timescale 1ns / 1ps
module full_adder(input a,input b,input cin,output sum,output cout);
    assign sum=a^b^cin;
    assign cout=(a&b)|(b&cin)|(cin&a);
endmodule
 
module main(input signed [9:0] A,B, output signed [19:0]product);
 wire [19:0]PP[0:9];
 wire [19:0]A_extended;
 wire [19:0]PP9_inverted;
 wire [19:0]sum_temp[0:8];
 wire cout_temp;
 
 assign A_extended={{10{A[9]}},A};
 
 genvar i;
 generate
 for(i=0;i<9;i=i+1) begin:pp_gen
 assign PP[i]=B[i]?(A_extended << i):20'b0;
 end
 endgenerate
 // Generate PP[9]
 assign PP[9]=A_extended << 9;
 // Invert PP[9] if B[9] is 1
 assign PP9_inverted = PP[9] ^ {20{B[9]}};
 // Sum all partial products using ripple carry adders
 rca_20 adder0(.a(PP[0]),.b(PP[1]),.cin(1'b0),.sum(sum_temp[0]),.cout(cout_temp));
 rca_20 adder1(.a(sum_temp[0]),.b(PP[2]),.cin(1'b0),.sum(sum_temp[1]),.cout(cout_temp));
 rca_20 adder2(.a(sum_temp[1]),.b(PP[3]),.cin(1'b0),.sum(sum_temp[2]),.cout(cout_temp));
 rca_20 adder3(.a(sum_temp[2]),.b(PP[4]),.cin(1'b0),.sum(sum_temp[3]),.cout(cout_temp));
 rca_20 adder4(.a(sum_temp[3]),.b(PP[5]),.cin(1'b0),.sum(sum_temp[4]),.cout(cout_temp));
 rca_20 adder5(.a(sum_temp[4]),.b(PP[6]),.cin(1'b0),.sum(sum_temp[5]),.cout(cout_temp));
 rca_20 adder6(.a(sum_temp[5]),.b(PP[7]),.cin(1'b0),.sum(sum_temp[6]),.cout(cout_temp));
 rca_20 adder7(.a(sum_temp[6]),.b(PP[8]),.cin(1'b0),.sum(sum_temp[7]),.cout(cout_temp));
 rca_20
adder8(.a(sum_temp[7]),.b(PP9_inverted),.cin(1'b0),.sum(sum_temp[8]),.cout(cout_temp));
 // Add B[9] as the carry-in for the final +1 adjustment
 rca_20 adder9(.a(sum_temp[8]),.b(20'b0),.cin(B[9]),.sum(product),.cout(cout_temp));
endmodule 

module rca_20(input [19:0] a,b,input cin,output[19:0]sum,output cout);
    wire [19:0] c;
    genvar i;
    generate
        for(i=0; i<20; i=i+1) begin: rca
            if(i==0)
                full_adder fa(.a(a[i]),.b(b[i]),.cin(cin),.sum(sum[i]),.cout(c[i]));
            else
                full_adder fa(.a(a[i]),.b(b[i]),.cin(c[i-1]),.sum(sum[i]),.cout(c[i]));
        end
    endgenerate
    assign cout=c[19];
endmodule